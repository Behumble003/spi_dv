//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
class spi_tlm extends uvm_sequence_item;

 `uvm_object_utils(spi_tlm)
 
  //
  // NEW
  //
  function new(string name = "spi_tlm");
    super.new(name);
  endfunction
  
endclass
